* NGSPICE file created from ShiftReg_row_10_2.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt TOP$1 VDD VSS Q PHI1 PHI2 D
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q PHI2 Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_1 D PHI1 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q VDD
+ VSS VDD VSS gf180mcu_fd_sc_mcu9t5v0__latq_1
.ends

.subckt ShiftReg_row_10_2 VDDd VSSd PHI_1 PHI_2 D_in Q[10] Q[4] Q[9] Q[3] Q[8] Q[5]
+ Q[7] Q[6] Q[2] Q[1]
XTOP$1_0[0] VDDd VSSd Q[1] PHI_1 PHI_2 D_in TOP$1
XTOP$1_0[1] VDDd VSSd Q[2] PHI_1 PHI_2 Q[1] TOP$1
XTOP$1_0[2] VDDd VSSd Q[3] PHI_1 PHI_2 Q[2] TOP$1
XTOP$1_0[3] VDDd VSSd Q[4] PHI_1 PHI_2 Q[3] TOP$1
XTOP$1_0[4] VDDd VSSd Q[5] PHI_1 PHI_2 Q[4] TOP$1
XTOP$1_0[5] VDDd VSSd Q[6] PHI_1 PHI_2 Q[5] TOP$1
XTOP$1_0[6] VDDd VSSd Q[7] PHI_1 PHI_2 Q[6] TOP$1
XTOP$1_0[7] VDDd VSSd Q[8] PHI_1 PHI_2 Q[7] TOP$1
XTOP$1_0[8] VDDd VSSd Q[9] PHI_1 PHI_2 Q[8] TOP$1
XTOP$1_0[9] VDDd VSSd Q[10] PHI_1 PHI_2 Q[9] TOP$1
.ends

