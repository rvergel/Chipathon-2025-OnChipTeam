** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/tb_swmatrix.sch
**.subckt tb_swmatrix
V1 VSSd GND 0
V2 VDDd VSSd {VDD}
xNO_ClkGen net2 clock_in net4 NO_ClkGen
x3 data datab VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x1 datab net6 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x4 clock clockb VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x5 clockb clock_in VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
xSWMATRIX data_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1] PIN[2] PIN[3]
+ PIN[4] PIN[5] PIN[6] PIN[7] PIN[8] PIN[9] PIN[10] PIN[11] PIN[12] PIN[13] PIN[14] PIN[15] PIN[16] PIN[17] PIN[18] PIN[19] PIN[20]
+ PIN[21] PIN[22] PIN[23] PIN[24] PIN[25] PIN[26] PIN[27] PIN[28] PIN[29] PIN[30] PIN[31] PIN[32] PIN[33] PIN[34] PIN[35] PIN[36] PIN[37]
+ PIN[38] PIN[39] PIN[40] PIN[41] PIN[42] PIN[43] PIN[44] PIN[45] PIN[46] PIN[47] PIN[48] swmatrix_48_by_10
* noconn D_out
* noconn BUS[1:10]
* noconn PIN[1:48]
x6 net2 net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x7 net1 PHI_2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x9 net4 net3 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x10 net3 PHI_1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x12 net6 net5 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x13 net5 data_in VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
**** begin user architecture code


.control

    save pin[1:48]
    TRAN 1n 100n
    write tb_swmatrix.raw

.endc



.include /foss/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/spice/gf180mcu_fd_sc_mcu9t5v0.spice
.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical



.param VDD = 1.8

.global VDDd VSSd

* clock
abit [ bit_node ]  input_vector
.model input_vector d_source(input_file="/foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/data_source/data_480.txt")
* data
aclock [ clock_node ] clock_vector
.model clock_vector d_source(input_file="/foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/data_source/data_480_clk.txt")
* convert digital signals to analog
aconvert [ bit_node clock_node ] [ data clock ] dac_in
.model dac_in dac_bridge (out_low=0V out_high=1.8V t_rise=0.2ns t_fall=0.2ns)


**** end user architecture code
**.ends

* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sym # of pins=3
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sch
.subckt NO_ClkGen PHI_2 CLK PHI_1
*.ipin CLK
*.opin PHI_2
*.opin PHI_1
x1 CLKB OUT_bot_d OUT_top VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
x2 OUT_top_d CLKbuf OUT_bot VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
x3 OUT_top PHI_2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x4 PHI_2 net3 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x5 net1 OUT_top_d VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x6 OUT_bot PHI_1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x7 PHI_1 net4 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x8 net2 OUT_bot_d VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x9 CLKB CLKbuf VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x10 CLK CLKB VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x11 net3 net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x12 net4 net2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_48_by_10/swmatrix_48_by_10.sym # of pins=6
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_48_by_10/swmatrix_48_by_10.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_48_by_10/swmatrix_48_by_10.sch
.subckt swmatrix_48_by_10 D_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1]
+ PIN[2] PIN[3] PIN[4] PIN[5] PIN[6] PIN[7] PIN[8] PIN[9] PIN[10] PIN[11] PIN[12] PIN[13] PIN[14] PIN[15] PIN[16] PIN[17] PIN[18] PIN[19]
+ PIN[20] PIN[21] PIN[22] PIN[23] PIN[24] PIN[25] PIN[26] PIN[27] PIN[28] PIN[29] PIN[30] PIN[31] PIN[32] PIN[33] PIN[34] PIN[35] PIN[36]
+ PIN[37] PIN[38] PIN[39] PIN[40] PIN[41] PIN[42] PIN[43] PIN[44] PIN[45] PIN[46] PIN[47] PIN[48]
*.iopin
*+ PIN[1],PIN[2],PIN[3],PIN[4],PIN[5],PIN[6],PIN[7],PIN[8],PIN[9],PIN[10],PIN[11],PIN[12],PIN[13],PIN[14],PIN[15],PIN[16],PIN[17],PIN[18],PIN[19],PIN[20],PIN[21],PIN[22],PIN[23],PIN[24],PIN[25],PIN[26],PIN[27],PIN[28],PIN[29],PIN[30],PIN[31],PIN[32],PIN[33],PIN[34],PIN[35],PIN[36],PIN[37],PIN[38],PIN[39],PIN[40],PIN[41],PIN[42],PIN[43],PIN[44],PIN[45],PIN[46],PIN[47],PIN[48]
*.iopin BUS[1],BUS[2],BUS[3],BUS[4],BUS[5],BUS[6],BUS[7],BUS[8],BUS[9],BUS[10]
*.ipin PHI_1
*.ipin PHI_2
*.ipin D_in
*.opin D_out
xswmatrix_row[1] D_in D_out_row[1] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1]
+ swmatrix_row_10
xswmatrix_row[2] D_out_row[1] D_out_row[2] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[2] swmatrix_row_10
xswmatrix_row[3] D_out_row[2] D_out_row[3] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[3] swmatrix_row_10
xswmatrix_row[4] D_out_row[3] D_out_row[4] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[4] swmatrix_row_10
xswmatrix_row[5] D_out_row[4] D_out_row[5] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[5] swmatrix_row_10
xswmatrix_row[6] D_out_row[5] D_out_row[6] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[6] swmatrix_row_10
xswmatrix_row[7] D_out_row[6] D_out_row[7] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[7] swmatrix_row_10
xswmatrix_row[8] D_out_row[7] D_out_row[8] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[8] swmatrix_row_10
xswmatrix_row[9] D_out_row[8] D_out_row[9] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[9] swmatrix_row_10
xswmatrix_row[10] D_out_row[9] D_out_row[10] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[10] swmatrix_row_10
xswmatrix_row[11] D_out_row[10] D_out_row[11] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[11] swmatrix_row_10
xswmatrix_row[12] D_out_row[11] D_out_row[12] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[12] swmatrix_row_10
xswmatrix_row[13] D_out_row[12] D_out_row[13] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[13] swmatrix_row_10
xswmatrix_row[14] D_out_row[13] D_out_row[14] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[14] swmatrix_row_10
xswmatrix_row[15] D_out_row[14] D_out_row[15] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[15] swmatrix_row_10
xswmatrix_row[16] D_out_row[15] D_out_row[16] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[16] swmatrix_row_10
xswmatrix_row[17] D_out_row[16] D_out_row[17] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[17] swmatrix_row_10
xswmatrix_row[18] D_out_row[17] D_out_row[18] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[18] swmatrix_row_10
xswmatrix_row[19] D_out_row[18] D_out_row[19] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[19] swmatrix_row_10
xswmatrix_row[20] D_out_row[19] D_out_row[20] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[20] swmatrix_row_10
xswmatrix_row[21] D_out_row[20] D_out_row[21] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[21] swmatrix_row_10
xswmatrix_row[22] D_out_row[21] D_out_row[22] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[22] swmatrix_row_10
xswmatrix_row[23] D_out_row[22] D_out_row[23] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[23] swmatrix_row_10
xswmatrix_row[24] D_out_row[23] D_out_row[24] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[24] swmatrix_row_10
xswmatrix_row[25] D_out_row[24] D_out_row[25] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[25] swmatrix_row_10
xswmatrix_row[26] D_out_row[25] D_out_row[26] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[26] swmatrix_row_10
xswmatrix_row[27] D_out_row[26] D_out_row[27] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[27] swmatrix_row_10
xswmatrix_row[28] D_out_row[27] D_out_row[28] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[28] swmatrix_row_10
xswmatrix_row[29] D_out_row[28] D_out_row[29] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[29] swmatrix_row_10
xswmatrix_row[30] D_out_row[29] D_out_row[30] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[30] swmatrix_row_10
xswmatrix_row[31] D_out_row[30] D_out_row[31] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[31] swmatrix_row_10
xswmatrix_row[32] D_out_row[31] D_out_row[32] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[32] swmatrix_row_10
xswmatrix_row[33] D_out_row[32] D_out_row[33] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[33] swmatrix_row_10
xswmatrix_row[34] D_out_row[33] D_out_row[34] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[34] swmatrix_row_10
xswmatrix_row[35] D_out_row[34] D_out_row[35] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[35] swmatrix_row_10
xswmatrix_row[36] D_out_row[35] D_out_row[36] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[36] swmatrix_row_10
xswmatrix_row[37] D_out_row[36] D_out_row[37] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[37] swmatrix_row_10
xswmatrix_row[38] D_out_row[37] D_out_row[38] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[38] swmatrix_row_10
xswmatrix_row[39] D_out_row[38] D_out_row[39] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[39] swmatrix_row_10
xswmatrix_row[40] D_out_row[39] D_out_row[40] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[40] swmatrix_row_10
xswmatrix_row[41] D_out_row[40] D_out_row[41] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[41] swmatrix_row_10
xswmatrix_row[42] D_out_row[41] D_out_row[42] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[42] swmatrix_row_10
xswmatrix_row[43] D_out_row[42] D_out_row[43] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[43] swmatrix_row_10
xswmatrix_row[44] D_out_row[43] D_out_row[44] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[44] swmatrix_row_10
xswmatrix_row[45] D_out_row[44] D_out_row[45] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[45] swmatrix_row_10
xswmatrix_row[46] D_out_row[45] D_out_row[46] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[46] swmatrix_row_10
xswmatrix_row[47] D_out_row[46] D_out_row[47] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[47] swmatrix_row_10
xswmatrix_row[48] D_out_row[47] D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[48]
+ swmatrix_row_10
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sym # of pins=6
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sch
.subckt swmatrix_row_10 D_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] pin
*.iopin pin
*.ipin PHI_2
*.ipin PHI_1
*.iopin BUS[1],BUS[2],BUS[3],BUS[4],BUS[5],BUS[6],BUS[7],BUS[8],BUS[9],BUS[10]
*.ipin D_in
*.opin D_out
xSR Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] D_out D_in PHI_1 PHI_2 ShiftReg_row_10_2
xTgates[1] Q[1] BUS[1] pin swmatrix_Tgate
xTgates[2] Q[2] BUS[2] pin swmatrix_Tgate
xTgates[3] Q[3] BUS[3] pin swmatrix_Tgate
xTgates[4] Q[4] BUS[4] pin swmatrix_Tgate
xTgates[5] Q[5] BUS[5] pin swmatrix_Tgate
xTgates[6] Q[6] BUS[6] pin swmatrix_Tgate
xTgates[7] Q[7] BUS[7] pin swmatrix_Tgate
xTgates[8] Q[8] BUS[8] pin swmatrix_Tgate
xTgates[9] Q[9] BUS[9] pin swmatrix_Tgate
xTgates[10] D_out BUS[10] pin swmatrix_Tgate
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sym # of pins=4
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sch
.subckt ShiftReg_row_10_2 Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] D_in PHI_1 PHI_2
*.ipin PHI_1
*.ipin PHI_2
*.ipin D_in
*.opin Q[1],Q[2],Q[3],Q[4],Q[5],Q[6],Q[7],Q[8],Q[9],Q[10]
xFF[1] D_in Q[1] PHI_1 PHI_2 DFF_2phase_1
xFF[2] Q[1] Q[2] PHI_1 PHI_2 DFF_2phase_1
xFF[3] Q[2] Q[3] PHI_1 PHI_2 DFF_2phase_1
xFF[4] Q[3] Q[4] PHI_1 PHI_2 DFF_2phase_1
xFF[5] Q[4] Q[5] PHI_1 PHI_2 DFF_2phase_1
xFF[6] Q[5] Q[6] PHI_1 PHI_2 DFF_2phase_1
xFF[7] Q[6] Q[7] PHI_1 PHI_2 DFF_2phase_1
xFF[8] Q[7] Q[8] PHI_1 PHI_2 DFF_2phase_1
xFF[9] Q[8] Q[9] PHI_1 PHI_2 DFF_2phase_1
xFF[10] Q[9] Q[10] PHI_1 PHI_2 DFF_2phase_1
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sym # of pins=3
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sch
.subckt swmatrix_Tgate control T2 T1
*.iopin T1
*.iopin T2
*.ipin control
* noconn control
* noconn T1
* noconn T2
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sym # of pins=4
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 D Q PHI_1 PHI_2
*.ipin D
*.ipin PHI_1
*.ipin PHI_2
*.opin Q
xmain D PHI_1 out_m VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
.ends

.GLOBAL GND
.end
