* Extracted by KLayout with GF180MCU LVS runset on : 11/08/2025 15:24

.SUBCKT ShiftReg_row_10_2 VSS D|Q D|Q|Q[2] D|Q|Q[3] D|Q|Q[4] D|Q|Q[5] D|Q|Q[9]
+ Q|Q[10] D|D_in E|PHI1 E|PHI2 D|Q|Q[1] D|Q|Q[6] D|Q|Q[7] D|Q|Q[8] VDD
M$1 VDD E|PHI1 \$2 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$2 \$3 \$2 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U PD=2.88U
M$3 VDD \$57 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$4 VDD E|PHI2 \$5 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$5 \$6 \$5 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U PD=2.88U
M$6 VDD \$60 D|Q|Q[1] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$7 VDD E|PHI1 \$7 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$8 \$8 \$7 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U PD=2.88U
M$9 VDD \$63 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$10 VDD E|PHI2 \$10 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$11 \$11 \$10 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$12 VDD \$65 D|Q|Q[2] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$13 VDD E|PHI1 \$13 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$14 \$14 \$13 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$15 VDD \$67 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$16 VDD E|PHI2 \$16 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$17 \$17 \$16 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$18 VDD \$69 D|Q|Q[3] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$19 VDD E|PHI1 \$19 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$20 \$20 \$19 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$21 VDD \$71 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$22 VDD E|PHI2 \$22 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$23 \$23 \$22 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$24 VDD \$73 D|Q|Q[4] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$25 VDD E|PHI1 \$25 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$26 \$26 \$25 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$27 VDD \$75 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$28 VDD E|PHI2 \$28 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$29 \$29 \$28 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$30 VDD \$77 D|Q|Q[5] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$31 VDD E|PHI1 \$31 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$32 \$32 \$31 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$33 VDD \$79 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$34 VDD E|PHI2 \$34 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$35 \$35 \$34 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$36 VDD \$81 D|Q|Q[6] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$37 VDD E|PHI1 \$36 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$38 \$37 \$36 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$39 VDD \$84 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$40 VDD E|PHI2 \$38 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$41 \$39 \$38 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$42 VDD \$87 D|Q|Q[7] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$43 VDD E|PHI1 \$40 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$44 \$41 \$40 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$45 VDD \$90 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$46 VDD E|PHI2 \$42 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$47 \$43 \$42 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$48 VDD \$93 D|Q|Q[8] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$49 VDD E|PHI1 \$44 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$50 \$45 \$44 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$51 VDD \$96 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$52 VDD E|PHI2 \$46 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$53 \$47 \$46 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$54 VDD \$99 D|Q|Q[9] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$55 VDD E|PHI1 \$49 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$56 \$50 \$49 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$57 VDD \$101 D|Q VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P PS=4.54U
+ PD=4.54U
M$58 VDD E|PHI2 \$52 VDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P PS=3.64U
+ PD=2.18U
M$59 \$53 \$52 VDD VDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$60 VDD \$103 Q|Q[10] VDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$61 \$238 D|D_in VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$62 \$57 \$2 \$238 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$63 \$57 \$3 \$240 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$64 VDD \$58 \$240 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$65 \$58 \$57 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$66 \$247 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$67 \$60 \$5 \$247 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$68 \$60 \$6 \$246 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$69 VDD \$61 \$246 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$70 \$61 \$60 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$71 \$255 D|Q|Q[1] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$72 \$63 \$7 \$255 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$73 \$63 \$8 \$254 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$74 VDD \$64 \$254 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$75 \$64 \$63 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$76 \$259 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$77 \$65 \$10 \$259 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$78 \$65 \$11 \$262 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$79 VDD \$66 \$262 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$80 \$66 \$65 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$81 \$267 D|Q|Q[2] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$82 \$67 \$13 \$267 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$83 \$67 \$14 \$270 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$84 VDD \$68 \$270 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$85 \$68 \$67 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$86 \$275 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$87 \$69 \$16 \$275 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$88 \$69 \$17 \$277 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$89 VDD \$70 \$277 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$90 \$70 \$69 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$91 \$284 D|Q|Q[3] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$92 \$71 \$19 \$284 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$93 \$71 \$20 \$285 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$94 VDD \$72 \$285 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$95 \$72 \$71 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$96 \$292 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U PD=1.24U
M$97 \$73 \$22 \$292 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$98 \$73 \$23 \$291 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$99 VDD \$74 \$291 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$100 \$74 \$73 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$101 \$297 D|Q|Q[4] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$102 \$75 \$25 \$297 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$103 \$75 \$26 \$300 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$104 VDD \$76 \$300 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$105 \$76 \$75 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$106 \$305 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$107 \$77 \$28 \$305 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$108 \$77 \$29 \$307 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$109 VDD \$78 \$307 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$110 \$78 \$77 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$111 \$312 D|Q|Q[5] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$112 \$79 \$31 \$312 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$113 \$79 \$32 \$315 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$114 VDD \$80 \$315 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$115 \$80 \$79 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$116 \$322 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$117 \$81 \$34 \$322 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$118 \$81 \$35 \$321 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$119 VDD \$82 \$321 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$120 \$82 \$81 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$121 \$327 D|Q|Q[6] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$122 \$84 \$36 \$327 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$123 \$84 \$37 \$330 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$124 VDD \$85 \$330 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$125 \$85 \$84 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$126 \$337 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$127 \$87 \$38 \$337 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$128 \$87 \$39 \$336 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$129 VDD \$88 \$336 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$130 \$88 \$87 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$131 \$342 D|Q|Q[7] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$132 \$90 \$40 \$342 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$133 \$90 \$41 \$345 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$134 VDD \$91 \$345 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$135 \$91 \$90 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$136 \$350 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$137 \$93 \$42 \$350 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$138 \$93 \$43 \$352 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$139 VDD \$94 \$352 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$140 \$94 \$93 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$141 \$359 D|Q|Q[8] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$142 \$96 \$44 \$359 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$143 \$96 \$45 \$360 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$144 VDD \$97 \$360 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P PS=2.08U
+ PD=1.9U
M$145 \$97 \$96 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$146 \$367 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$147 \$99 \$46 \$367 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$148 \$99 \$47 \$366 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$149 VDD \$100 \$366 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$150 \$100 \$99 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P PS=1.9U
+ PD=3.64U
M$151 \$375 D|Q|Q[9] VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$152 \$101 \$49 \$375 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$153 \$101 \$50 \$374 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$154 VDD \$102 \$374 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$155 \$102 \$101 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$156 \$381 D|Q VDD VDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$157 \$103 \$52 \$381 VDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$158 \$103 \$53 \$382 VDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$159 VDD \$104 \$382 VDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$160 \$104 \$103 VDD VDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$161 VSS \$57 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$162 VSS \$60 D|Q|Q[1] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$163 VSS \$63 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$164 VSS \$65 D|Q|Q[2] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$165 VSS \$67 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$166 VSS \$69 D|Q|Q[3] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$167 VSS \$71 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$168 VSS \$73 D|Q|Q[4] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$169 VSS \$75 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$170 VSS \$77 D|Q|Q[5] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$171 VSS \$79 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$172 VSS \$81 D|Q|Q[6] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$173 VSS \$84 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$174 VSS \$87 D|Q|Q[7] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$175 VSS \$90 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$176 VSS \$93 D|Q|Q[8] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$177 VSS \$96 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$178 VSS \$99 D|Q|Q[9] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$179 VSS \$101 D|Q VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P PS=3.52U
+ PD=3.52U
M$180 VSS \$103 Q|Q[10] VSS nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$181 VSS E|PHI1 \$2 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P PS=2.46U
+ PD=1.49U
M$182 \$3 \$2 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$183 VSS E|PHI2 \$5 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P PS=2.46U
+ PD=1.49U
M$184 \$6 \$5 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$185 VSS E|PHI1 \$7 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P PS=2.46U
+ PD=1.49U
M$186 \$8 \$7 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$187 VSS E|PHI2 \$10 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$188 \$11 \$10 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$189 VSS E|PHI1 \$13 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$190 \$14 \$13 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$191 VSS E|PHI2 \$16 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$192 \$17 \$16 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$193 VSS E|PHI1 \$19 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$194 \$20 \$19 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$195 VSS E|PHI2 \$22 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$196 \$23 \$22 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$197 VSS E|PHI1 \$25 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$198 \$26 \$25 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$199 VSS E|PHI2 \$28 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$200 \$29 \$28 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$201 VSS E|PHI1 \$31 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$202 \$32 \$31 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$203 VSS E|PHI2 \$34 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$204 \$35 \$34 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$205 VSS E|PHI1 \$36 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$206 \$37 \$36 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$207 VSS E|PHI2 \$38 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$208 \$39 \$38 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$209 VSS E|PHI1 \$40 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$210 \$41 \$40 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$211 VSS E|PHI2 \$42 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$212 \$43 \$42 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$213 VSS E|PHI1 \$44 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$214 \$45 \$44 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$215 VSS E|PHI2 \$46 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$216 \$47 \$46 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$217 VSS E|PHI1 \$49 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$218 \$50 \$49 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$219 VSS E|PHI2 \$52 VSS nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$220 \$53 \$52 VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$221 \$108 D|D_in VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$222 \$57 \$3 \$108 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$223 \$109 \$2 \$57 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$224 VSS \$58 \$109 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$225 \$58 \$57 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$226 \$117 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$227 \$60 \$6 \$117 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$228 \$116 \$5 \$60 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$229 VSS \$61 \$116 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$230 \$61 \$60 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$231 \$125 D|Q|Q[1] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$232 \$63 \$8 \$125 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$233 \$126 \$7 \$63 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$234 VSS \$64 \$126 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$235 \$64 \$63 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$236 \$133 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$237 \$65 \$11 \$133 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$238 \$132 \$10 \$65 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$239 VSS \$66 \$132 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$240 \$66 \$65 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$241 \$144 D|Q|Q[2] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$242 \$67 \$14 \$144 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$243 \$145 \$13 \$67 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$244 VSS \$68 \$145 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$245 \$68 \$67 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$246 \$150 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$247 \$69 \$17 \$150 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$248 \$152 \$16 \$69 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$249 VSS \$70 \$152 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$250 \$70 \$69 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$251 \$160 D|Q|Q[3] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$252 \$71 \$20 \$160 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$253 \$161 \$19 \$71 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$254 VSS \$72 \$161 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$255 \$72 \$71 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$256 \$167 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$257 \$73 \$23 \$167 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$258 \$168 \$22 \$73 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$259 VSS \$74 \$168 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$260 \$74 \$73 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$261 \$177 D|Q|Q[4] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$262 \$75 \$26 \$177 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$263 \$178 \$25 \$75 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$264 VSS \$76 \$178 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$265 \$76 \$75 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$266 \$186 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$267 \$77 \$29 \$186 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$268 \$184 \$28 \$77 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$269 VSS \$78 \$184 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$270 \$78 \$77 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$271 \$195 D|Q|Q[5] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$272 \$79 \$32 \$195 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$273 \$197 \$31 \$79 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$274 VSS \$80 \$197 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$275 \$80 \$79 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$276 \$202 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$277 \$81 \$35 \$202 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$278 \$203 \$34 \$81 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$279 VSS \$82 \$203 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$280 \$82 \$81 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$281 \$211 D|Q|Q[6] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$282 \$84 \$37 \$211 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$283 \$214 \$36 \$84 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$284 VSS \$85 \$214 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$285 \$85 \$84 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$286 \$220 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$287 \$87 \$39 \$220 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$288 \$219 \$38 \$87 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$289 VSS \$88 \$219 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$290 \$88 \$87 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$291 \$230 D|Q|Q[7] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$292 \$90 \$41 \$230 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$293 \$229 \$40 \$90 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$294 VSS \$91 \$229 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$295 \$91 \$90 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$296 \$227 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$297 \$93 \$43 \$227 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$298 \$223 \$42 \$93 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$299 VSS \$94 \$223 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$300 \$94 \$93 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$301 \$196 D|Q|Q[8] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$302 \$96 \$45 \$196 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$303 \$194 \$44 \$96 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$304 VSS \$97 \$194 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P PS=1.49U
+ PD=1.31U
M$305 \$97 \$96 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P PS=1.31U
+ PD=2.46U
M$306 \$171 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$307 \$99 \$47 \$171 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$308 \$175 \$46 \$99 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$309 VSS \$100 \$175 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$310 \$100 \$99 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$311 \$143 D|Q|Q[9] VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$312 \$101 \$50 \$143 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$313 \$142 \$49 \$101 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$314 VSS \$102 \$142 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$315 \$102 \$101 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$316 \$122 D|Q VSS VSS nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$317 \$103 \$53 \$122 VSS nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$318 \$118 \$52 \$103 VSS nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$319 VSS \$104 \$118 VSS nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$320 \$104 \$103 VSS VSS nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
.ENDS ShiftReg_row_10_2
