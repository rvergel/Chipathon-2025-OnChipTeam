** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/tb_swmatrix.sch
**.subckt tb_swmatrix
Vvssd VSSd GND 0
Vvddd VDDd VSSd {VDD}
xNO_ClkGen net9 net10 net11 net12 net13 NO_ClkGen
x3 data datab VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x1 datab net6 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x4 clock clockb VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
x5 clockb clock_in VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_2
xSWMATRIX data_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1] PIN[2] PIN[3]
+ PIN[4] PIN[5] VDDd VSSd enable swmatrix_5_by_10
* noconn D_out
* noconn BUS[1:10]
* noconn PIN[1:5]
x6 net2 net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x7 net1 PHI_2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x9 net4 net3 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x10 net3 PHI_1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x12 net6 net5 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x13 net5 data_in VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
x2 net8 net7 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_4
x8 net7 enable VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_8
Venable net8 VSSd 0
**** begin user architecture code


.control

    save all
    TRAN 0.2n 350n
    write tb_swmatrix.raw

.endc



.include /foss/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/spice/gf180mcu_fd_sc_mcu9t5v0.spice
.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical



.param VDD = 3.3

*.global VDDd VSSd

* clock
abit [ bit_node ]  input_vector
.model input_vector d_source(input_file="/foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/data_source/data_swmatrix5_10.txt")
* data
aclock [ clock_node ] clock_vector
.model clock_vector d_source(input_file="/foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/testbenches/data_source/data_swmatrix5_10_clk.txt")
* convert digital signals to analog
aconvert [ bit_node clock_node ] [ data clock ] dac_in
.model dac_in dac_bridge (out_low=0V out_high=3.3V t_rise=0.2ns t_fall=0.2ns)


**** end user architecture code
**.ends

* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sym # of pins=5
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/NO_ClkGen/NO_ClkGen.sch
.subckt NO_ClkGen PHI_2 CLK PHI_1 VDDd VSSd
*.ipin CLK
*.opin PHI_2
*.opin PHI_1
*.iopin VDDd
*.iopin VSSd
x1 CLKB OUT_bot_d OUT_top VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
x2 OUT_top_d CLKbuf OUT_bot VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
x3 OUT_top PHI_2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x4 PHI_2 net5 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x5 net3 net2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x6 OUT_bot PHI_1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x7 PHI_1 net6 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x8 net4 net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x9 CLKB CLKbuf VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x10 CLK CLKB VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x11 net5 net3 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x12 net6 net4 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x13 net2 net7 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x15 net1 net8 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x17 net7 net9 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x18 net8 net12 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x14 net9 net10 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x16 net12 net11 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x19 net10 OUT_top_d VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x20 net11 OUT_bot_d VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
* noconn VDDd
* noconn VSSd
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_5_by_10/swmatrix_5_by_10.sym # of pins=9
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_5_by_10/swmatrix_5_by_10.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_5_by_10/swmatrix_5_by_10.sch
.subckt swmatrix_5_by_10 D_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1]
+ PIN[2] PIN[3] PIN[4] PIN[5] VDDd VSSd enable
*.iopin PIN[1],PIN[2],PIN[3],PIN[4],PIN[5]
*.iopin BUS[1],BUS[2],BUS[3],BUS[4],BUS[5],BUS[6],BUS[7],BUS[8],BUS[9],BUS[10]
*.ipin PHI_1
*.ipin PHI_2
*.ipin D_in
*.opin D_out
*.iopin VDDd
*.iopin VSSd
*.ipin enable
xswmatrix_row[1] D_in D_out_row[1] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[1] VDDd
+ VSSd enable swmatrix_row_10
xswmatrix_row[2] D_out_row[1] D_out_row[2] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[2] VDDd VSSd enable swmatrix_row_10
xswmatrix_row[3] D_out_row[2] D_out_row[3] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[3] VDDd VSSd enable swmatrix_row_10
xswmatrix_row[4] D_out_row[3] D_out_row[4] PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10]
+ PIN[4] VDDd VSSd enable swmatrix_row_10
xswmatrix_row[5] D_out_row[4] D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] PIN[5] VDDd
+ VSSd enable swmatrix_row_10
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sym # of pins=9
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_row_10/swmatrix_row_10.sch
.subckt swmatrix_row_10 D_in D_out PHI_1 PHI_2 BUS[1] BUS[2] BUS[3] BUS[4] BUS[5] BUS[6] BUS[7] BUS[8] BUS[9] BUS[10] pin VDDd
+ VSSd enable
*.iopin pin
*.ipin PHI_2
*.ipin PHI_1
*.iopin BUS[1],BUS[2],BUS[3],BUS[4],BUS[5],BUS[6],BUS[7],BUS[8],BUS[9],BUS[10]
*.ipin D_in
*.opin D_out
*.iopin VDDd
*.iopin VSSd
*.ipin enable
xSR Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] D_out D_in PHI_1 PHI_2 VDDd VSSd ShiftReg_row_10_2
xTgates[1] Q[1] BUS[1] pin VDDd VSSd enable swmatrix_Tgate
xTgates[2] Q[2] BUS[2] pin VDDd VSSd enable swmatrix_Tgate
xTgates[3] Q[3] BUS[3] pin VDDd VSSd enable swmatrix_Tgate
xTgates[4] Q[4] BUS[4] pin VDDd VSSd enable swmatrix_Tgate
xTgates[5] Q[5] BUS[5] pin VDDd VSSd enable swmatrix_Tgate
xTgates[6] Q[6] BUS[6] pin VDDd VSSd enable swmatrix_Tgate
xTgates[7] Q[7] BUS[7] pin VDDd VSSd enable swmatrix_Tgate
xTgates[8] Q[8] BUS[8] pin VDDd VSSd enable swmatrix_Tgate
xTgates[9] Q[9] BUS[9] pin VDDd VSSd enable swmatrix_Tgate
xTgates[10] D_out BUS[10] pin VDDd VSSd enable swmatrix_Tgate
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sym # of pins=6
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/ShiftReg_row_10_2/ShiftReg_row_10_2.sch
.subckt ShiftReg_row_10_2 Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] Q[9] Q[10] D_in PHI_1 PHI_2 VDDd VSSd
*.ipin PHI_1
*.ipin PHI_2
*.ipin D_in
*.opin Q[1],Q[2],Q[3],Q[4],Q[5],Q[6],Q[7],Q[8],Q[9],Q[10]
*.iopin VDDd
*.iopin VSSd
xFF[1] D_in Q[1] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[2] Q[1] Q[2] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[3] Q[2] Q[3] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[4] Q[3] Q[4] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[5] Q[4] Q[5] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[6] Q[5] Q[6] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[7] Q[6] Q[7] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[8] Q[7] Q[8] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[9] Q[8] Q[9] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
xFF[10] Q[9] Q[10] PHI_1 PHI_2 VDDd VSSd DFF_2phase_1
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sym # of pins=6
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/swmatrix_Tgate/swmatrix_Tgate.sch
.subckt swmatrix_Tgate control T2 T1 VDDd VSSd enable
*.iopin T1
*.iopin T2
*.iopin VDDd
*.iopin VSSd
*.ipin control
*.ipin enable
XM1 T1 gated_control T2 VSSd nfet_03v3 L=0.28u W=mn_w nf=6 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 T1 gated_controlb T2 VDDd pfet_03v3 L=0.28u W=mp_w nf=6 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
**** begin user architecture code


.param mn_w=24u
.param mp_w=72u

**** end user architecture code
x1 gated_control gated_controlb VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
x2 control enable net1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__nand2_1
x3 net1 gated_control VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
.ends


* expanding   symbol:  Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sym # of pins=6
** sym_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/Chipathon-2025-OnChipTeam/designs/switch_matrix/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 D Q PHI_1 PHI_2 VDDd VSSd
*.ipin D
*.ipin PHI_1
*.ipin PHI_2
*.opin Q
*.iopin VDDd
*.iopin VSSd
xmain D PHI_1 out_m VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
* noconn VSSd
* noconn VDDd
.ends

.GLOBAL GND
.end
